V1 1 0 5
R1 1 2 1K
R2 2 3 2K
R3 3 0 3K
.DC V1 6 6 1
.PRINT DC V1(2,3) V(2) I(R2)
.END